library verilog;
use verilog.vl_types.all;
entity MIPS is
    port(
        clk             : in     vl_logic;
        nrst            : in     vl_logic
    );
end MIPS;
